version https://git-lfs.github.com/spec/v1
oid sha256:725453c493a2c5a781bf0540776478203838a607dee6dfc475166d60ce22750d
size 13731
