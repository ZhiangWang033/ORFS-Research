version https://git-lfs.github.com/spec/v1
oid sha256:59ec3093031fcea1808cc8bd8f3dfeef120b49343a626e016791d7dad0e23f24
size 2460509
