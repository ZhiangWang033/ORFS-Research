version https://git-lfs.github.com/spec/v1
oid sha256:5a30e0626b465841101b96edba94e3b7c145fb0c5d3bc5bd7efc55ce1cac6a1a
size 14058
