version https://git-lfs.github.com/spec/v1
oid sha256:14337b02358a90f84d9f4844bc8ea3778459a1bf145c5e7fe6a9583467edc79f
size 24467
